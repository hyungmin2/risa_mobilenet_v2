`ifndef __DEFINES_VH__
`define __DEFINES_VH__

`define CEILDIV(x,y) (((x) + (y) -1)/(y))
`define MAX(x,y) ( ( (x) > (y) ) ? (x) : (y) )
`define MIN(x,y) ( ( (x) < (y) ) ? (x) : (y) )

 
`endif //__DEFINES_VH__